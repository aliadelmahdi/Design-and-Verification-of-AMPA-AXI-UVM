package AXI_env_pkg;

    import  uvm_pkg::*;
    import shared_pkg::*;

    `include "AXI_config.sv"
    `include "AXI_master_pkg.sv"
    `include "AXI_slave_pkg.sv"
    `include "AXI_coverage_collector.sv"
    `include "AXI_scoreboard.sv"
    `include "AXI_env.sv"

endpackage : AXI_env_pkg