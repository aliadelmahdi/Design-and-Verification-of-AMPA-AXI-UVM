package AXI_env_pkg;

    import  uvm_pkg::*;
    import shared_pkg::*;

    `include "AXI_config.svh"
    `include "AXI_master_pkg.svh"
    `include "AXI_slave_pkg.svh"
    `include "AXI_coverage_collector.svh"
    `include "AXI_scoreboard.svh"
    `include "AXI_env.svh"

endpackage : AXI_env_pkg