`ifndef AXI_MASTER_PKG_SVH
`define AXI_MASTER_PKG_SVH

    `include "AXI_master_seq_item.svh"
    `include "AXI_master_sequences.svh"
    `include "AXI_master_driver.svh"
    `include "AXI_master_monitor.svh"
    `include "AXI_master_sequencer.svh"
    `include "AXI_master_agent.svh"

`endif // AXI_MASTER_PKG_SVH