`include "axi_defines.svh" // For macros
import shared_pkg::*; // For enums and parameters

module golden_model ();

endmodule : golden_model
