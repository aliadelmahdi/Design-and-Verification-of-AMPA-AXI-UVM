import shared_pkg::*; // For enums and parameters

`include "AXI_master_gld.sv"
`include "AXI_slave_gld.sv"