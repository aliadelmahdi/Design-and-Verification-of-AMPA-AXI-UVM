`ifndef AXI_MASTER_SEQUENCES_SV
`define AXI_MASTER_SEQUENCES_SV

    `include "AXI_master_reset_sequence.sv"
    `include "AXI_master_main_sequence.sv"

`endif // AXI_MASTER_SEQUENCES_SV
