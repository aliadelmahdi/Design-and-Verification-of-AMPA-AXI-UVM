// The following `define` values represent bit widths and sizes used in the design. 
// are only for convenience and to make the code more readable. 
import shared_pkg::*; // For enums and parameters

`include "AXI_master.sv"
`include "AXI_slave.sv"