`ifndef AXI_SLAVE_SEQUENCES_SVH
`define AXI_SLAVE_SEQUENCES_SVH

    `include "AXI_slave_main_sequence.svh"

`endif // AXI_SLAVE_SEQUENCES_SVH