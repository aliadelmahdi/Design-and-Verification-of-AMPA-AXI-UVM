
package AXI_test_pkg;

    import  uvm_pkg::*;
    import  shared_pkg::*;
    import  AXI_env_pkg::*;
    
    `include "AXI_test_base.sv"

endpackage : AXI_test_pkg