`ifndef AXI_MASTER_SEQUENCES_SVH
`define AXI_MASTER_SEQUENCES_SVH

    `include "AXI_master_reset_sequence.svh"
    `include "AXI_master_main_sequence.svh"

`endif // AXI_MASTER_SEQUENCES_SVH
