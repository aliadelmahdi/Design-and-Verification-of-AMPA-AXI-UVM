`ifndef AXI_SLAVE_SV
`define AXI_SLAVE_SV

module AXI_slave ();

endmodule

`endif // AXI_SLAVE_SV