import shared_pkg::*; // For enums and parameters

`include "AXI_master.sv"
`include "AXI_slave.sv"