`ifndef AXI_SLAVE_SEQUENCES_SV
`define AXI_SLAVE_SEQUENCES_SV

    `include "AXI_slave_main_sequence.sv"

`endif // AXI_SLAVE_SEQUENCES_SV