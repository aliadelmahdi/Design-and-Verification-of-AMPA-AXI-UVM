// ============================================================================
// Read-after-write (RAW) sequence
// ============================================================================
`ifndef AXI_MASTER_READ_AFTER_WRITE_SEQ_SVH
`define AXI_MASTER_READ_AFTER_WRITE_SEQ_SVH

// Writes to an address range, then reads it back to check coherency.
class AXI_master_read_after_write_seq extends AXI_master_main_sequence;

    `uvm_object_utils(AXI_master_read_after_write_seq)

    function new(string name = "AXI_master_read_after_write_seq");
        super.new(name);
    endfunction : new

    task body;
        repeat(`TEST_ITER_SMALL) begin
            // Phase 1: WRITE
            configure_seq_item();
            start_item(seq_item);
            // TODO: write phase constraints
            // assert(seq_item.randomize() with { is_write == 1; }) else ...
            assert(seq_item.randomize()) else $error("Master Randomization Failed");
            finish_item(seq_item);

            // Phase 2: READ (same region)
            configure_seq_item();
            start_item(seq_item);
            // TODO: make read target the same address window as write
            // assert(seq_item.randomize() with { is_read == 1; same_region_as_prev == 1; }) else ...
            assert(seq_item.randomize()) else $error("Master Randomization Failed");
            finish_item(seq_item);
        end
    endtask : body

endclass : AXI_master_read_after_write_seq

`endif // AXI_MASTER_READ_AFTER_WRITE_SEQ_SVH