`ifndef AXI_SLAVE_SEQUENCES_SVH
`define AXI_SLAVE_SEQUENCES_SVH

// AXI Slave Sequences Package - includes all predefined slave sequences
`include "AXI_slave_main_sequence.svh" // Main randomized slave response sequence

`endif // AXI_SLAVE_SEQUENCES_SVH
