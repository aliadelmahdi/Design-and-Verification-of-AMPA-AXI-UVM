package AXI_test_pkg;

    // Import required packages
    import uvm_pkg::*;      // UVM base classes and utilities
    import shared_pkg::*;   // Shared typedefs, parameters, and constants
    import AXI_env_pkg::*;  // AXI environment and its components
    
    // Include test files
    `include "AXI_test_base.svh" // Base AXI test definition

endpackage : AXI_test_pkg