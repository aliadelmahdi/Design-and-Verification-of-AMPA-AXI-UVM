// ============================================================================
// Write-after-read (WAR) sequence
// ============================================================================
`ifndef AXI_MASTER_WRITE_AFTER_READ_SEQ_SVH
`define AXI_MASTER_WRITE_AFTER_READ_SEQ_SVH

// Reads a region, then writes to it (ordering/latency interaction).
class AXI_master_write_after_read_seq extends AXI_master_main_sequence;

    `uvm_object_utils(AXI_master_write_after_read_seq)

    function new(string name = "AXI_master_write_after_read_seq");
        super.new(name);
    endfunction : new

    task body;
        repeat(`TEST_ITER_SMALL) begin
            // Phase 1: READ
            configure_seq_item();
            start_item(seq_item);
            // TODO: read constraints
            // assert(seq_item.randomize() with { is_read == 1; }) else ...
            assert(seq_item.randomize()) else $error("Master Randomization Failed");
            finish_item(seq_item);

            // Phase 2: WRITE (same/overlapping region)
            configure_seq_item();
            start_item(seq_item);
            // TODO: write to same/overlapping region
            // assert(seq_item.randomize() with { is_write == 1; same_region_as_prev == 1; }) else ...
            assert(seq_item.randomize()) else $error("Master Randomization Failed");
            finish_item(seq_item);
        end
    endtask : body

endclass : AXI_master_write_after_read_seq

`endif // AXI_MASTER_WRITE_AFTER_READ_SEQ_SVH