`ifndef AXI_MASTER_PKG_SV
`define AXI_MASTER_PKG_SV

    `include "AXI_master_seq_item.sv"
    `include "AXI_master_sequences.sv"
    `include "AXI_master_driver.sv"
    `include "AXI_master_monitor.sv"
    `include "AXI_master_sequencer.sv"
    `include "AXI_master_agent.sv"

`endif // AXI_MASTER_PKG_SV